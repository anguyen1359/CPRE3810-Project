library ieee;
use ieee.std_logic_1164.all;

entity decoder5to32 is
  port (
    i_D : in  std_logic_vector(4 downto 0);  -- 5-bit input
    o_Q : out std_logic_vector(31 downto 0)  -- 32-bit one-hot output
  );
end entity decoder5to32;

architecture dataflow of decoder5to32 is
begin
  with i_D select
    o_Q <= "00000000000000000000000000000001" when "00000", -- 0
           "00000000000000000000000000000010" when "00001", -- 1
           "00000000000000000000000000000100" when "00010", -- 2
           "00000000000000000000000000001000" when "00011", -- 3
           "00000000000000000000000000010000" when "00100", -- 4
	   "00000000000000000000000000100000" when "00101", -- 5
           "00000000000000000000000001000000" when "00110", -- 6
           "00000000000000000000000010000000" when "00111", -- 7
           "00000000000000000000000100000000" when "01000", -- 8
           "00000000000000000000001000000000" when "01001", -- 9
	   "00000000000000000000010000000000" when "01010", -- 10
           "00000000000000000000100000000000" when "01011", -- 11
           "00000000000000000001000000000000" when "01100", -- 12
           "00000000000000000010000000000000" when "01101", -- 13
           "00000000000000000100000000000000" when "01110", -- 14
	   "00000000000000001000000000000000" when "01111", -- 15
           "00000000000000010000000000000000" when "10000", -- 16
           "00000000000000100000000000000000" when "10001", -- 17
           "00000000000001000000000000000000" when "10010", -- 18
           "00000000000010000000000000000000" when "10011", -- 19
	   "00000000000100000000000000000000" when "10100", -- 20
           "00000000001000000000000000000000" when "10101", -- 21
           "00000000010000000000000000000000" when "10110", -- 22
           "00000000100000000000000000000000" when "10111", -- 23
           "00000001000000000000000000000000" when "11000", -- 24
	   "00000010000000000000000000000000" when "11001", -- 25
           "00000100000000000000000000000000" when "11010", -- 26
           "00001000000000000000000000000000" when "11011", -- 27
           "00010000000000000000000000000000" when "11100", -- 28
           "00100000000000000000000000000000" when "11101", -- 29
	   "01000000000000000000000000000000" when "11110", -- 30      
           "10000000000000000000000000000000" when "11111", -- 31
           (others => '0') when others; -- default
end architecture dataflow;

